parameter R_TYPE    = 3'b000;
parameter I_TYPE    = 3'b001;
parameter L_TYPE    = 3'b010;
parameter S_TYPE    = 3'b011;
parameter B_TYPE    = 3'b100;
parameter J_TYPE    = 3'b101;
parameter U_TYPE    = 3'b101;
parameter MATH_TYPE = 3'b101;
parameter BM_TYPE   = 3'b101;
parameter M_TYPE    = 3'b110;
