module mem_manage(mem_r, mem_w, addr, )